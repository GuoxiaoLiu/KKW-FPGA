library ieee;
use ieee.std_logic_1164.all;
library work;
use work.lowmc_pkg.all;

package debug_pkg is
    -- lowmc parameter
    constant PL : std_logic_vector(N - 1 downto 0) := "010101010101010101010100000001010001000001000101000001010101010100000100010001010101010100010001000000000001000100000100000100010";
    constant CI : std_logic_vector(N - 1 downto 0) := "010101010101010101010100000001010001000001000101000001010101010100000100010001010101010100010001000000000001000100000100000100010";
    constant KE : std_logic_vector(N - 1 downto 0) := "010101010101010101010100000001010001000001000101000001010101010100000100010001010101010100010001000000000001000100000100000100010";
    constant ME : std_logic_vector(512 - 1 downto 0) := "00000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001000000010000000100000001";
    
    
    
end debug_pkg;
